module main;
  initial
    begin
      $display("Hello, World!");
      $finish(0);
    end
endmodule
