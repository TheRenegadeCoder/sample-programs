module main

fn main(){
	println('Hello, world!')
}